`include "design.v"

module AWMC_tb();
    reg clk, reset, start, pause,lid;
    wire [2:0] stage;
    wire done;
    wire lido;

    AWMC uut(.clk(clk),.reset(reset),.start(start),.pause(pause),.stage(stage),.done(done),.lid(lid));

    initial begin
        reset = 1'b0;
        #1
        reset = 1'b1;
        #1
        reset = 1'b0;
        clk = 1'b0;

        forever #5 clk = ~clk;
    end

    initial begin
        start = 1'b0;
        pause = 1'b0;

        $dumpfile("tb.vcd");
        $dumpvars(0,AWMC_tb);

        #10
        start = 1'b1;
        lid = 1'b1;
        #20
        start = 1'b0;
        #100
        pause = 1'b1;
        lid = 1'b0;
        #105
        pause = 1'b0;
        #110
        start = 1'b0;
        #120 
        start = 1'b0;
        #150
        reset = 1'b0;
        #155
        start = 1'b0;
        lid = 1'b1;
        #160
        start = 1'b0;
        #165
        lid = 1'b1;
        #167
        lid = 1'b0;
        #170
        pause = 1'b0;
        #200
        reset = 1'b1;
        start = 1'b1;
        lid = 1'b1;
        #205
        reset = 1'b0;  
        #240
        start = 1'b0;
        lid = 1'b0;
        #250
        pause = 1'b1;
        #310
        pause = 1'b0;
        lid = 1'b1;
        #360
        lid = 1'b0;

        #400 $finish;

    end

endmodule
